//axi 3
`define FIXED    2'b00
`define INCR     2'b01
`define WRAP     2'b10
`define REVERSE  2'b11

`define OKAY     2'b00
`define EXOKAY   2'b01
`define SLVERR   2'b10
`define DECERR   2'b11

`define SLV0_START_ADDR 0
`define SLV0_END_ADDR 4095
`define SLV1_START_ADDR 4096
`define SLV1_END_ADDR 8191
`define SLV2_START_ADDR 8192
`define SLV2_END_ADDR 12287
`define SLV3_START_ADDR 12288
`define SLV3_END_ADDR 16383

`define SLV0 2'b01
`define SLV1 2'b10
`define SLV2 2'b11

`define MST0 2'b01
`define MST1 2'b10
`define MST2 2'b11

//ahb
`define IDLE    2'b00
`define BUSY    2'b01
`define NONSEQ  2'b10
`define SEQ     2'b11